`ifndef _MPCACHE_H_
`define _MPCACHE_H_

`define IN_PORT_NUM         (16)
`define OUT_PORT_NUM        (16)
`define DATA_WIDTH          (32)
    
`define DA_WIDTH            (4)
`define PRORITY_WIDTH       (3)
`define BLK_ADDR_WIDTH      (14)
`define BLK_R_TIMES_WIDTH   (4)
`define BLK_W_TIMES_WIDTH   (4)

`endif