`ifndef _MPCACHE_H_
`define _MPCACHE_H_

`define IN_PORT_NUM         (16)
`define OUT_PORT_NUM        (16)
`define DATA_WIDTH          (32)
    
`define DA_WIDTH            (4)
`define PRORITY_WIDTH       (3)
`define BLK_ADDR_WIDTH      (10)

`endif